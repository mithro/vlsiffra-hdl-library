/**
Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

     http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
 */

/** DO NOT EDIT -- This file is generated by `make_techmap_v.py` file **/

(* techmap_celltype = "$add" *)
module _map_add(A, B, Y);

    parameter A_SIGNED = 0;
    parameter B_SIGNED = 0;
    parameter A_WIDTH = 1;
    parameter B_WIDTH = 1;
    parameter Y_WIDTH = 1;

    (* force_downto *)
    input [A_WIDTH-1:0] A;
    (* force_downto *)
    input [B_WIDTH-1:0] B;
    (* force_downto *)
    output [Y_WIDTH-1:0] Y;

    // Simple sanity checks
    //wire _TECHMAP_FAIL_ = A_WIDTH != Y_WIDTH;
    //wire _TECHMAP_FAIL_ = B_WIDTH != Y_WIDTH;

    genvar i;
    generate
        if (A_WIDTH == 2)
            add_b02 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 3)
            add_b03 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 4)
            add_b04 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 5)
            add_b05 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 6)
            add_b06 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 7)
            add_b07 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 8)
            add_b08 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 9)
            add_b09 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 10)
            add_b10 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 11)
            add_b11 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 12)
            add_b12 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 13)
            add_b13 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 14)
            add_b14 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 15)
            add_b15 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 16)
            add_b16 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 17)
            add_b17 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 18)
            add_b18 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 19)
            add_b19 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 20)
            add_b20 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 21)
            add_b21 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 22)
            add_b22 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 23)
            add_b23 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 24)
            add_b24 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 25)
            add_b25 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 26)
            add_b26 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 27)
            add_b27 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 28)
            add_b28 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 29)
            add_b29 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 30)
            add_b30 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 31)
            add_b31 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 32)
            add_b32 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 33)
            add_b33 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 34)
            add_b34 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 35)
            add_b35 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 36)
            add_b36 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 37)
            add_b37 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 38)
            add_b38 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 39)
            add_b39 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 40)
            add_b40 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 41)
            add_b41 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 42)
            add_b42 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 43)
            add_b43 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 44)
            add_b44 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 45)
            add_b45 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 46)
            add_b46 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 47)
            add_b47 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 48)
            add_b48 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 49)
            add_b49 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 50)
            add_b50 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 51)
            add_b51 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 52)
            add_b52 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 53)
            add_b53 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 54)
            add_b54 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 55)
            add_b55 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 56)
            add_b56 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 57)
            add_b57 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 58)
            add_b58 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 59)
            add_b59 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 60)
            add_b60 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 61)
            add_b61 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 62)
            add_b62 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
        else if (A_WIDTH == 63)
            add_b63 _TECHMAP_REPLACE_ (.a(A), .b(B), .o(Y));
    endgenerate
endmodule
