/* 2-bit wide adder */
(* blackbox *)
module add_b02(
	input [1:0] a,
	input [1:0] b,
	output [1:0] o);
endmodule

/* 3-bit wide adder */
(* blackbox *)
module add_b03(
	input [2:0] a,
	input [2:0] b,
	output [2:0] o);
endmodule

/* 4-bit wide adder */
(* blackbox *)
module add_b04(
	input [3:0] a,
	input [3:0] b,
	output [3:0] o);
endmodule

/* 5-bit wide adder */
(* blackbox *)
module add_b05(
	input [4:0] a,
	input [4:0] b,
	output [4:0] o);
endmodule

/* 6-bit wide adder */
(* blackbox *)
module add_b06(
	input [5:0] a,
	input [5:0] b,
	output [5:0] o);
endmodule

/* 7-bit wide adder */
(* blackbox *)
module add_b07(
	input [6:0] a,
	input [6:0] b,
	output [6:0] o);
endmodule

/* 8-bit wide adder */
(* blackbox *)
module add_b08(
	input [7:0] a,
	input [7:0] b,
	output [7:0] o);
endmodule

/* 9-bit wide adder */
(* blackbox *)
module add_b09(
	input [8:0] a,
	input [8:0] b,
	output [8:0] o);
endmodule

/* 10-bit wide adder */
(* blackbox *)
module add_b10(
	input [9:0] a,
	input [9:0] b,
	output [9:0] o);
endmodule

/* 11-bit wide adder */
(* blackbox *)
module add_b11(
	input [10:0] a,
	input [10:0] b,
	output [10:0] o);
endmodule

/* 12-bit wide adder */
(* blackbox *)
module add_b12(
	input [11:0] a,
	input [11:0] b,
	output [11:0] o);
endmodule

/* 13-bit wide adder */
(* blackbox *)
module add_b13(
	input [12:0] a,
	input [12:0] b,
	output [12:0] o);
endmodule

/* 14-bit wide adder */
(* blackbox *)
module add_b14(
	input [13:0] a,
	input [13:0] b,
	output [13:0] o);
endmodule

/* 15-bit wide adder */
(* blackbox *)
module add_b15(
	input [14:0] a,
	input [14:0] b,
	output [14:0] o);
endmodule

/* 16-bit wide adder */
(* blackbox *)
module add_b16(
	input [15:0] a,
	input [15:0] b,
	output [15:0] o);
endmodule

/* 17-bit wide adder */
(* blackbox *)
module add_b17(
	input [16:0] a,
	input [16:0] b,
	output [16:0] o);
endmodule

/* 18-bit wide adder */
(* blackbox *)
module add_b18(
	input [17:0] a,
	input [17:0] b,
	output [17:0] o);
endmodule

/* 19-bit wide adder */
(* blackbox *)
module add_b19(
	input [18:0] a,
	input [18:0] b,
	output [18:0] o);
endmodule

/* 20-bit wide adder */
(* blackbox *)
module add_b20(
	input [9:0] a,
	input [9:0] b,
	output [9:0] o);
endmodule

/* 21-bit wide adder */
(* blackbox *)
module add_b21(
	input [20:0] a,
	input [20:0] b,
	output [20:0] o);
endmodule

/* 22-bit wide adder */
(* blackbox *)
module add_b22(
	input [21:0] a,
	input [21:0] b,
	output [21:0] o);
endmodule

/* 23-bit wide adder */
(* blackbox *)
module add_b23(
	input [22:0] a,
	input [22:0] b,
	output [22:0] o);
endmodule

/* 24-bit wide adder */
(* blackbox *)
module add_b24(
	input [23:0] a,
	input [23:0] b,
	output [23:0] o);
endmodule

/* 25-bit wide adder */
(* blackbox *)
module add_b25(
	input [24:0] a,
	input [24:0] b,
	output [24:0] o);
endmodule

/* 26-bit wide adder */
(* blackbox *)
module add_b26(
	input [25:0] a,
	input [25:0] b,
	output [25:0] o);
endmodule

/* 27-bit wide adder */
(* blackbox *)
module add_b27(
	input [26:0] a,
	input [26:0] b,
	output [26:0] o);
endmodule

/* 28-bit wide adder */
(* blackbox *)
module add_b28(
	input [27:0] a,
	input [27:0] b,
	output [27:0] o);
endmodule

/* 29-bit wide adder */
(* blackbox *)
module add_b29(
	input [28:0] a,
	input [28:0] b,
	output [28:0] o);
endmodule
