(* blackbox *)
module add_b02(
	input [1:0] a,
	input [1:0] b,
	output [1:0] o);
endmodule

(* blackbox *)
module add_b03(
	input [2:0] a,
	input [2:0] b,
	output [2:0] o);
endmodule

(* blackbox *)
module add_b04(
	input [3:0] a,
	input [3:0] b,
	output [3:0] o);
endmodule

(* blackbox *)
module add_b05(
	input [4:0] a,
	input [4:0] b,
	output [4:0] o);
endmodule

(* blackbox *)
module add_b06(
	input [5:0] a,
	input [5:0] b,
	output [5:0] o);
endmodule

(* blackbox *)
module add_b07(
	input [6:0] a,
	input [6:0] b,
	output [6:0] o);
endmodule

(* blackbox *)
module add_b08(
	input [7:0] a,
	input [7:0] b,
	output [7:0] o);
endmodule

(* blackbox *)
module add_b09(
	input [8:0] a,
	input [8:0] b,
	output [8:0] o);
endmodule

(* blackbox *)
module add_b10(
	input [9:0] a,
	input [9:0] b,
	output [9:0] o);
endmodule

(* blackbox *)
module add_b11(
	input [10:0] a,
	input [10:0] b,
	output [10:0] o);
endmodule

(* blackbox *)
module add_b12(
	input [11:0] a,
	input [11:0] b,
	output [11:0] o);
endmodule

(* blackbox *)
module add_b13(
	input [12:0] a,
	input [12:0] b,
	output [12:0] o);
endmodule

(* blackbox *)
module add_b14(
	input [13:0] a,
	input [13:0] b,
	output [13:0] o);
endmodule

(* blackbox *)
module add_b15(
	input [14:0] a,
	input [14:0] b,
	output [14:0] o);
endmodule

(* blackbox *)
module add_b16(
	input [15:0] a,
	input [15:0] b,
	output [15:0] o);
endmodule

(* blackbox *)
module add_b17(
	input [16:0] a,
	input [16:0] b,
	output [16:0] o);
endmodule

(* blackbox *)
module add_b18(
	input [17:0] a,
	input [17:0] b,
	output [17:0] o);
endmodule

(* blackbox *)
module add_b19(
	input [18:0] a,
	input [18:0] b,
	output [18:0] o);
endmodule
