/**
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *      http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

/** DO NOT EDIT -- This file is generated by `make_bb_v.py` file **/


/* 2-bit wide adder */
(* blackbox *)
module add_b02 (
        input [2:0] a,
        input [2:0] b,
        output [2:0] o);
endmodule

/* 3-bit wide adder */
(* blackbox *)
module add_b03 (
        input [3:0] a,
        input [3:0] b,
        output [3:0] o);
endmodule

/* 4-bit wide adder */
(* blackbox *)
module add_b04 (
        input [4:0] a,
        input [4:0] b,
        output [4:0] o);
endmodule

/* 5-bit wide adder */
(* blackbox *)
module add_b05 (
        input [5:0] a,
        input [5:0] b,
        output [5:0] o);
endmodule

/* 6-bit wide adder */
(* blackbox *)
module add_b06 (
        input [6:0] a,
        input [6:0] b,
        output [6:0] o);
endmodule

/* 7-bit wide adder */
(* blackbox *)
module add_b07 (
        input [7:0] a,
        input [7:0] b,
        output [7:0] o);
endmodule

/* 8-bit wide adder */
(* blackbox *)
module add_b08 (
        input [8:0] a,
        input [8:0] b,
        output [8:0] o);
endmodule

/* 9-bit wide adder */
(* blackbox *)
module add_b09 (
        input [9:0] a,
        input [9:0] b,
        output [9:0] o);
endmodule

/* 10-bit wide adder */
(* blackbox *)
module add_b10 (
        input [10:0] a,
        input [10:0] b,
        output [10:0] o);
endmodule

/* 11-bit wide adder */
(* blackbox *)
module add_b11 (
        input [11:0] a,
        input [11:0] b,
        output [11:0] o);
endmodule

/* 12-bit wide adder */
(* blackbox *)
module add_b12 (
        input [12:0] a,
        input [12:0] b,
        output [12:0] o);
endmodule

/* 13-bit wide adder */
(* blackbox *)
module add_b13 (
        input [13:0] a,
        input [13:0] b,
        output [13:0] o);
endmodule

/* 14-bit wide adder */
(* blackbox *)
module add_b14 (
        input [14:0] a,
        input [14:0] b,
        output [14:0] o);
endmodule

/* 15-bit wide adder */
(* blackbox *)
module add_b15 (
        input [15:0] a,
        input [15:0] b,
        output [15:0] o);
endmodule

/* 16-bit wide adder */
(* blackbox *)
module add_b16 (
        input [16:0] a,
        input [16:0] b,
        output [16:0] o);
endmodule

/* 17-bit wide adder */
(* blackbox *)
module add_b17 (
        input [17:0] a,
        input [17:0] b,
        output [17:0] o);
endmodule

/* 18-bit wide adder */
(* blackbox *)
module add_b18 (
        input [18:0] a,
        input [18:0] b,
        output [18:0] o);
endmodule

/* 19-bit wide adder */
(* blackbox *)
module add_b19 (
        input [19:0] a,
        input [19:0] b,
        output [19:0] o);
endmodule

/* 20-bit wide adder */
(* blackbox *)
module add_b20 (
        input [20:0] a,
        input [20:0] b,
        output [20:0] o);
endmodule

/* 21-bit wide adder */
(* blackbox *)
module add_b21 (
        input [21:0] a,
        input [21:0] b,
        output [21:0] o);
endmodule

/* 22-bit wide adder */
(* blackbox *)
module add_b22 (
        input [22:0] a,
        input [22:0] b,
        output [22:0] o);
endmodule

/* 23-bit wide adder */
(* blackbox *)
module add_b23 (
        input [23:0] a,
        input [23:0] b,
        output [23:0] o);
endmodule

/* 24-bit wide adder */
(* blackbox *)
module add_b24 (
        input [24:0] a,
        input [24:0] b,
        output [24:0] o);
endmodule

/* 25-bit wide adder */
(* blackbox *)
module add_b25 (
        input [25:0] a,
        input [25:0] b,
        output [25:0] o);
endmodule

/* 26-bit wide adder */
(* blackbox *)
module add_b26 (
        input [26:0] a,
        input [26:0] b,
        output [26:0] o);
endmodule

/* 27-bit wide adder */
(* blackbox *)
module add_b27 (
        input [27:0] a,
        input [27:0] b,
        output [27:0] o);
endmodule

/* 28-bit wide adder */
(* blackbox *)
module add_b28 (
        input [28:0] a,
        input [28:0] b,
        output [28:0] o);
endmodule

/* 29-bit wide adder */
(* blackbox *)
module add_b29 (
        input [29:0] a,
        input [29:0] b,
        output [29:0] o);
endmodule

/* 30-bit wide adder */
(* blackbox *)
module add_b30 (
        input [30:0] a,
        input [30:0] b,
        output [30:0] o);
endmodule

/* 31-bit wide adder */
(* blackbox *)
module add_b31 (
        input [31:0] a,
        input [31:0] b,
        output [31:0] o);
endmodule

/* 32-bit wide adder */
(* blackbox *)
module add_b32 (
        input [32:0] a,
        input [32:0] b,
        output [32:0] o);
endmodule

/* 33-bit wide adder */
(* blackbox *)
module add_b33 (
        input [33:0] a,
        input [33:0] b,
        output [33:0] o);
endmodule

/* 34-bit wide adder */
(* blackbox *)
module add_b34 (
        input [34:0] a,
        input [34:0] b,
        output [34:0] o);
endmodule

/* 35-bit wide adder */
(* blackbox *)
module add_b35 (
        input [35:0] a,
        input [35:0] b,
        output [35:0] o);
endmodule

/* 36-bit wide adder */
(* blackbox *)
module add_b36 (
        input [36:0] a,
        input [36:0] b,
        output [36:0] o);
endmodule

/* 37-bit wide adder */
(* blackbox *)
module add_b37 (
        input [37:0] a,
        input [37:0] b,
        output [37:0] o);
endmodule

/* 38-bit wide adder */
(* blackbox *)
module add_b38 (
        input [38:0] a,
        input [38:0] b,
        output [38:0] o);
endmodule

/* 39-bit wide adder */
(* blackbox *)
module add_b39 (
        input [39:0] a,
        input [39:0] b,
        output [39:0] o);
endmodule

/* 40-bit wide adder */
(* blackbox *)
module add_b40 (
        input [40:0] a,
        input [40:0] b,
        output [40:0] o);
endmodule

/* 41-bit wide adder */
(* blackbox *)
module add_b41 (
        input [41:0] a,
        input [41:0] b,
        output [41:0] o);
endmodule

/* 42-bit wide adder */
(* blackbox *)
module add_b42 (
        input [42:0] a,
        input [42:0] b,
        output [42:0] o);
endmodule

/* 43-bit wide adder */
(* blackbox *)
module add_b43 (
        input [43:0] a,
        input [43:0] b,
        output [43:0] o);
endmodule

/* 44-bit wide adder */
(* blackbox *)
module add_b44 (
        input [44:0] a,
        input [44:0] b,
        output [44:0] o);
endmodule

/* 45-bit wide adder */
(* blackbox *)
module add_b45 (
        input [45:0] a,
        input [45:0] b,
        output [45:0] o);
endmodule

/* 46-bit wide adder */
(* blackbox *)
module add_b46 (
        input [46:0] a,
        input [46:0] b,
        output [46:0] o);
endmodule

/* 47-bit wide adder */
(* blackbox *)
module add_b47 (
        input [47:0] a,
        input [47:0] b,
        output [47:0] o);
endmodule

/* 48-bit wide adder */
(* blackbox *)
module add_b48 (
        input [48:0] a,
        input [48:0] b,
        output [48:0] o);
endmodule

/* 49-bit wide adder */
(* blackbox *)
module add_b49 (
        input [49:0] a,
        input [49:0] b,
        output [49:0] o);
endmodule

/* 50-bit wide adder */
(* blackbox *)
module add_b50 (
        input [50:0] a,
        input [50:0] b,
        output [50:0] o);
endmodule

/* 51-bit wide adder */
(* blackbox *)
module add_b51 (
        input [51:0] a,
        input [51:0] b,
        output [51:0] o);
endmodule

/* 52-bit wide adder */
(* blackbox *)
module add_b52 (
        input [52:0] a,
        input [52:0] b,
        output [52:0] o);
endmodule

/* 53-bit wide adder */
(* blackbox *)
module add_b53 (
        input [53:0] a,
        input [53:0] b,
        output [53:0] o);
endmodule

/* 54-bit wide adder */
(* blackbox *)
module add_b54 (
        input [54:0] a,
        input [54:0] b,
        output [54:0] o);
endmodule

/* 55-bit wide adder */
(* blackbox *)
module add_b55 (
        input [55:0] a,
        input [55:0] b,
        output [55:0] o);
endmodule

/* 56-bit wide adder */
(* blackbox *)
module add_b56 (
        input [56:0] a,
        input [56:0] b,
        output [56:0] o);
endmodule

/* 57-bit wide adder */
(* blackbox *)
module add_b57 (
        input [57:0] a,
        input [57:0] b,
        output [57:0] o);
endmodule

/* 58-bit wide adder */
(* blackbox *)
module add_b58 (
        input [58:0] a,
        input [58:0] b,
        output [58:0] o);
endmodule

/* 59-bit wide adder */
(* blackbox *)
module add_b59 (
        input [59:0] a,
        input [59:0] b,
        output [59:0] o);
endmodule

/* 60-bit wide adder */
(* blackbox *)
module add_b60 (
        input [60:0] a,
        input [60:0] b,
        output [60:0] o);
endmodule

/* 61-bit wide adder */
(* blackbox *)
module add_b61 (
        input [61:0] a,
        input [61:0] b,
        output [61:0] o);
endmodule

/* 62-bit wide adder */
(* blackbox *)
module add_b62 (
        input [62:0] a,
        input [62:0] b,
        output [62:0] o);
endmodule

/* 63-bit wide adder */
(* blackbox *)
module add_b63 (
        input [63:0] a,
        input [63:0] b,
        output [63:0] o);
endmodule
